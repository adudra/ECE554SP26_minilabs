module fifo_tb();

// SIGNAL DECLARATION //
logic clk;
logic rst_n;
logic rden;
logic wren;
logic [7:0] i_data;
logic [7:0] o_data;
logic full;
logic empty;

// DUT INSTANTIATION //
FIFO #(.DEPTH(8), .DATA_WIDTH(8)) 
    ififo(
    .clk(clk),
    .rst_n(rst_n), 
    .rden(rden),
    .wren(wren),
    .i_data(i_data),
    .o_data(o_data),
    .full(full),
    .empty(empty)
);

// STIMULUS APPLICATION //
initial begin
    // INITIAL CONDITIONS //
    clk = 1'b0;
    rst_n = 1'b0;
    rden = 1'b0;
    wren = 1'b0;
    i_data = 1'b0;

    // TEST BEGIN BELOW //
    @(negedge clk) begin 
	rst_n = 1'b1; //de-assert reset 
	i_data = 8'h11;
    end 

    // CASE 1: enables held low, data inputted (no data written, and empty flag high
    @(posedge clk) 
    if (o_data !== 6'h00) begin 
	$disply("FAILURE CASE1: outputted content was non-zero upon reset");
	$stop();
    end 
    if (!empty) begin 
	$disply("FAILURE CASE1: empty flag did not assert when fifo was empty");
	$stop();
    end

    // CASE 2: write enable high, read enable low 
    @(negedge clk) wren = 1'b1;

    @(posedge clk);
    #1
    if (ififo.fifo_mem[0] !== 8'h11) begin 
	$display("FAILURE CASE2: did not correctly write data to fifo when wren enabled");
	$stop();
    end 

    // CASE 3: write enable low, read enable high 
    @(negedge clk) begin 
	wren = 1'b0;
	rden = 1'b1;
    end

    @(posedge clk);
    #1
    if (o_data !== 8'h11) begin 
	$display("FAILURE CASE3: did not correctly read data from fifo");
	$stop();
    end 
    if (!empty) begin 
	$display("FAILURE CASE3: did not correctly detect empty fifo");
	$stop();
    end 

    // CASE 4: write enable high, read enable high
    @(negedge clk) begin 
	wren = 1'b1;
        rden = 1'b0; //deasserting rden to fill fifo buffer
        i_data = 8'h22;
    end

    repeat (3) @(posedge clk); //fill fifo buffer with 3 instances of 8'h22

    @(negedge clk) begin 
	rden = 1'b1;
    end

    @(posedge clk);
    #1 
    if (o_data !== 8'h22) begin 
	$display("FAILURE CASE4: did not correctly read data from fifo when both enables asserted");
	$stop();
    end
    if (ififo.w_ptr !== 3'h5) begin //internal check to confirm correctly read and wrote simultaneously
	$display("FAILURE CASE4: write pointer was not expected when both enables asserted");
	$stop();
    end
    if (ififo.r_ptr !== 3'h2) begin //internal check to confirm correctly read and wrote simultaneously 
	$display("FAILURE CASE4: read pointer was not expected when both enables asserted");
	$stop();
    end

   // CASE 5: ensure full flag correctly sets
   @(negedge clk) begin 
	rden = 1'b0;
	i_data = 8'h33;
   end 

   repeat (5) @(posedge clk);

   #1 
   if (!full) begin 
	$display("FAILURE CASE5: full flag not asserted when fifo should be full");
	$stop();
   end 

   $display("YAHOO! All tests passed");
   $stop();
end

// CLOCK GENERATION //
always begin
 #5 clk <= ~clk;
end

endmodule