module baud_rate_generator(
    input clk,
    input rst,
    output tx_en,
    output rx_en,
    output reg [15:0] baud_divisor
);



endmodule