module convolution_tb();
    
endmodule